module decoder4to16 (w, y);
    input [3:0] w;
    output [15:0] y;
    reg [15:0] y;
    always @(*)
    begin
        case(w)
            0: y = 16'b0000000000000001;
            1: y = 16'b0000000000000010;
            2: y = 16'b0000000000000100;
            3: y = 16'b0000000000001000;
            4: y = 16'b0000000000010000;
            5: y = 16'b0000000000100000;
            6: y = 16'b0000000001000000;
            7: y = 16'b0000000010000000;
            8: y = 16'b0000000100000000;
            9: y = 16'b0000001000000000;
            10: y = 16'b0000010000000000;
            11: y = 16'b0000100000000000;
            12: y = 16'b0001000000000000;
            13: y = 16'b0010000000000000;
            14: y = 16'b0100000000000000;
            15: y = 16'b1000000000000000;
        endcase
    end
endmodule