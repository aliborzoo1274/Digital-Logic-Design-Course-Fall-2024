`timescale 1ns/1ns
module Top_Module_Tb ();
    reg [15:0] inp1, inp2;
    reg [2:0] opc;
    wire [15:0] out;
    wire overflow;
    Top_Module UT (inp1, inp2, opc, out, overflow);
    initial
    begin
        inp1 = 16'b0000000000000100;
        inp2 = 16'b0000000000001000;
        opc = 3'b001;
        #5;

        inp1 = 16'b0000000000100000;
        inp2 = 16'b0000000000010000;
        opc = 3'b001;
        #5;

        inp1 = 16'b0000000010000000;
        inp2 = 16'b0000000000000100;
        opc = 3'b010;
        #5;

        inp1 = 16'b1000000000000000;
        inp2 = 16'b0000000010000000;
        opc = 3'b010;
        #5;

        inp1 = 16'b0000000001000000;
        inp2 = 16'b0000000000000001;
        opc = 3'b011;
        #5;

        inp1 = 16'b0010000000000000;
        inp2 = 16'b0100000000000000;
        opc = 3'b011;
        #5;

        inp1 = 16'b0000000000000000;
        inp2 = 16'b0000000000010000;
        opc = 3'b100;
        #5;

        inp1 = 16'b0000000000010000;
        inp2 = 16'b0000100000000000;
        opc = 3'b100;
        #5;

        inp1 = 16'b0000000000001000;
        inp2 = 16'b1000000000000000;
        opc = 3'b101;
        #5;

        inp1 = 16'b0000000001000000;
        inp2 = 16'b1000000000000000;
        opc = 3'b101;
        #5;

        inp1 = 16'b0000000000000010;
        inp2 = 16'b0010000000000000;
        opc = 3'b110;
        #5;

        inp1 = 16'b0000000000010000;
        inp2 = 16'b0000000000100000;
        opc = 3'b110;
        #5;

        inp1 = 16'b0000000010000000;
        inp2 = 16'b0000001000000000;
        opc = 3'b111;
        #5;

        inp1 = 16'b0000000000000000;
        inp2 = 16'b0100000000000000;
        opc = 3'b111;
        #5;
    end
endmodule